module controlUnit(
    input wire clk,
    input wire reset,
)

endmodule