module cpu(
    input wire clk, reset
);

    //single bit wires
    wire PCWrite;
    wire PCWriteCond;
    wire EPCWrite;
    wire MultDiv;

    // TO DO
    // 1. Add the mux control signals
    


endmodule