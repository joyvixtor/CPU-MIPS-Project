module controlUnit(
    input wire clk,
    input wire reset,

    //STATES
    parameter ST_ADD = 6'b000000, //0
    parameter ST_ADDI = 6'b000001, //1
)

endmodule